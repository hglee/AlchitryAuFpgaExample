/**
 * @file fifo.sv
 * @brief Top level FIFO module
 *
 * Origin from FPGA Prototyping by SystemVerilog Examples - Pong P. Chu
 */
`begin_keywords "1800-2017"
`timescale 1ns/1ps

module fifo
  #(
    parameter DATA_WIDTH = 8, // number of bits in a word
    ADDR_WIDTH = 4 // number of address bits
    )
   (
    input logic                   clk, reset,
    input logic                   rd, wr,
    input logic [DATA_WIDTH-1:0]  w_data,
    output logic                  empty, full,
    output logic [DATA_WIDTH-1:0] r_data
    );

   // signal
   logic [ADDR_WIDTH-1:0]         w_addr, r_addr;
   logic                          wr_en, full_tmp;

   // body
   // write enabled only when FIFO is not full
   assign wr_en = wr & ~full_tmp;
   assign full = full_tmp;

   // instantiate fifo control unit
   fifo_ctrl #(.ADDR_WIDTH(ADDR_WIDTH)) c_unit (.*, .full(full_tmp));

   // instantiate register file
   reg_file #(.DATA_WIDTH(DATA_WIDTH), .ADDR_WIDTH(ADDR_WIDTH)) f_unit (.*);

endmodule: fifo

`end_keywords
