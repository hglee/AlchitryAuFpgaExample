/**
 * @file top.sv
 * @brief top level without FIFO HDL
 */
module top
  (
   input logic clk,
   input logic rst_n,
   output logic [7:0] led,
   input logic ft_clk,
   input logic ft_rxf_n, // rx full
   input logic ft_txe_n, // tx empty
   output logic [15:0] ft_data, // data
   output logic [1:0] ft_be,  // byte enable
   output logic ft_rd_n, // read enable
   output logic ft_wr_n, // write enable
   output logic ft_oe_n // output enable
   );

   logic [15:0] din_reg, din_next;
   logic        wr_reg, wr_next;
   logic [7:0]  led_reg, led_next;

   always_ff @(posedge ft_clk)
     begin
        if (rst_n)
          begin
             // not reset
             din_reg <= din_next;
             wr_reg <= wr_next;
             led_reg <= led_next;
          end
        else
          begin
             // reset
             din_reg <= 0;
             wr_reg <= 0;
             led_reg <= 0;
          end
     end

   always_comb
     begin
        if (ft_txe_n)
          begin
             din_next = din_reg;
             wr_next = 1;
             led_next = 8'h01;
          end
        else
          begin
             // increase if empty
             din_next = din_reg + 1;
             wr_next = 0;
             led_next = 8'hf1;
          end
     end

   // output
   assign led = led_reg;
   assign ft_data = din_reg;
   assign ft_be = 2'b11;
   assign ft_rd_n = 1;
   assign ft_wr_n = wr_reg;
   assign ft_oe_n = 1;

endmodule // top
